// Copyright 2021 The CFU-Playground Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.



module Cfu (
  input               cmd_valid,
  output              cmd_ready,
  input      [9:0]    cmd_payload_function_id,
  input      [31:0]   cmd_payload_inputs_0,
  input      [31:0]   cmd_payload_inputs_1,
  output reg          rsp_valid,
  input               rsp_ready,
  output reg [31:0]   rsp_payload_outputs_0,
  input               reset,
  input               clk
);

  reg [31:0] EXP_LOOKUP_TABLE [0:511];

  initial begin
      EXP_LOOKUP_TABLE[0] = 32'h7fffffff;
      EXP_LOOKUP_TABLE[1] = 32'h7C0FD5AA;
      EXP_LOOKUP_TABLE[2] = 32'h783EAFEF;
      EXP_LOOKUP_TABLE[3] = 32'h748B9A80;
      EXP_LOOKUP_TABLE[4] = 32'h70F5A893;
      EXP_LOOKUP_TABLE[5] = 32'h6D7BF4A7;
      EXP_LOOKUP_TABLE[6] = 32'h6A1DA04B;
      EXP_LOOKUP_TABLE[7] = 32'h66D9D3E3;
      EXP_LOOKUP_TABLE[8] = 32'h63AFBE7A;
      EXP_LOOKUP_TABLE[9] = 32'h609E9586;
      EXP_LOOKUP_TABLE[10] = 32'h5DA594B7;
      EXP_LOOKUP_TABLE[11] = 32'h5AC3FDCB;
      EXP_LOOKUP_TABLE[12] = 32'h57F91857;
      EXP_LOOKUP_TABLE[13] = 32'h5544319F;
      EXP_LOOKUP_TABLE[14] = 32'h52A49C64;
      EXP_LOOKUP_TABLE[15] = 32'h5019B0BF;
      EXP_LOOKUP_TABLE[16] = 32'h4DA2CBF1;
      EXP_LOOKUP_TABLE[17] = 32'h4B3F503E;
      EXP_LOOKUP_TABLE[18] = 32'h48EEA4C3;
      EXP_LOOKUP_TABLE[19] = 32'h46B03552;
      EXP_LOOKUP_TABLE[20] = 32'h4483724D;
      EXP_LOOKUP_TABLE[21] = 32'h4267D07F;
      EXP_LOOKUP_TABLE[22] = 32'h405CC8FF;
      EXP_LOOKUP_TABLE[23] = 32'h3E61D906;
      EXP_LOOKUP_TABLE[24] = 32'h3C7681D7;
      EXP_LOOKUP_TABLE[25] = 32'h3A9A4899;
      EXP_LOOKUP_TABLE[26] = 32'h38CCB63C;
      EXP_LOOKUP_TABLE[27] = 32'h370D5757;
      EXP_LOOKUP_TABLE[28] = 32'h355BBC12;
      EXP_LOOKUP_TABLE[29] = 32'h33B77803;
      EXP_LOOKUP_TABLE[30] = 32'h32202217;
      EXP_LOOKUP_TABLE[31] = 32'h30955477;
      EXP_LOOKUP_TABLE[32] = 32'h2F16AC6C;
      EXP_LOOKUP_TABLE[33] = 32'h2DA3CA4B;
      EXP_LOOKUP_TABLE[34] = 32'h2C3C515A;
      EXP_LOOKUP_TABLE[35] = 32'h2ADFE7B7;
      EXP_LOOKUP_TABLE[36] = 32'h298E3648;
      EXP_LOOKUP_TABLE[37] = 32'h2846E89E;
      EXP_LOOKUP_TABLE[38] = 32'h2709ACE4;
      EXP_LOOKUP_TABLE[39] = 32'h25D633C9;
      EXP_LOOKUP_TABLE[40] = 32'h24AC306E;
      EXP_LOOKUP_TABLE[41] = 32'h238B584F;
      EXP_LOOKUP_TABLE[42] = 32'h22736336;
      EXP_LOOKUP_TABLE[43] = 32'h21640B24;
      EXP_LOOKUP_TABLE[44] = 32'h205D0C41;
      EXP_LOOKUP_TABLE[45] = 32'h1F5E24CC;
      EXP_LOOKUP_TABLE[46] = 32'h1E67150B;
      EXP_LOOKUP_TABLE[47] = 32'h1D779F37;
      EXP_LOOKUP_TABLE[48] = 32'h1C8F8772;
      EXP_LOOKUP_TABLE[49] = 32'h1BAE93B5;
      EXP_LOOKUP_TABLE[50] = 32'h1AD48BC2;
      EXP_LOOKUP_TABLE[51] = 32'h1A013915;
      EXP_LOOKUP_TABLE[52] = 32'h193466DA;
      EXP_LOOKUP_TABLE[53] = 32'h186DE1DA;
      EXP_LOOKUP_TABLE[54] = 32'h17AD7873;
      EXP_LOOKUP_TABLE[55] = 32'h16F2FA8A;
      EXP_LOOKUP_TABLE[56] = 32'h163E397E;
      EXP_LOOKUP_TABLE[57] = 32'h158F081D;
      EXP_LOOKUP_TABLE[58] = 32'h14E53A9C;
      EXP_LOOKUP_TABLE[59] = 32'h1440A685;
      EXP_LOOKUP_TABLE[60] = 32'h13A122B3;
      EXP_LOOKUP_TABLE[61] = 32'h13068744;
      EXP_LOOKUP_TABLE[62] = 32'h1270AD90;
      EXP_LOOKUP_TABLE[63] = 32'h11DF7020;
      EXP_LOOKUP_TABLE[64] = 32'h1152AAA3;
      EXP_LOOKUP_TABLE[65] = 32'h10CA39E9;
      EXP_LOOKUP_TABLE[66] = 32'h1045FBD3;
      EXP_LOOKUP_TABLE[67] = 32'h0FC5CF52;
      EXP_LOOKUP_TABLE[68] = 32'h0F49945A;
      EXP_LOOKUP_TABLE[69] = 32'h0ED12BDB;
      EXP_LOOKUP_TABLE[70] = 32'h0E5C77BB;
      EXP_LOOKUP_TABLE[71] = 32'h0DEB5ACC;
      EXP_LOOKUP_TABLE[72] = 32'h0D7DB8C7;
      EXP_LOOKUP_TABLE[73] = 32'h0D137641;
      EXP_LOOKUP_TABLE[74] = 32'h0CAC78AB;
      EXP_LOOKUP_TABLE[75] = 32'h0C48A644;
      EXP_LOOKUP_TABLE[76] = 32'h0BE7E616;
      EXP_LOOKUP_TABLE[77] = 32'h0B8A1FF2;
      EXP_LOOKUP_TABLE[78] = 32'h0B2F3C65;
      EXP_LOOKUP_TABLE[79] = 32'h0AD724B7;
      EXP_LOOKUP_TABLE[80] = 32'h0A81C2E0;
      EXP_LOOKUP_TABLE[81] = 32'h0A2F0188;
      EXP_LOOKUP_TABLE[82] = 32'h09DECBFD;
      EXP_LOOKUP_TABLE[83] = 32'h09910E33;
      EXP_LOOKUP_TABLE[84] = 32'h0945B4B9;
      EXP_LOOKUP_TABLE[85] = 32'h08FCACB9;
      EXP_LOOKUP_TABLE[86] = 32'h08B5E3F0;
      EXP_LOOKUP_TABLE[87] = 32'h087148AB;
      EXP_LOOKUP_TABLE[88] = 32'h082EC9C4;
      EXP_LOOKUP_TABLE[89] = 32'h07EE569A;
      EXP_LOOKUP_TABLE[90] = 32'h07AFDF11;
      EXP_LOOKUP_TABLE[91] = 32'h07735389;
      EXP_LOOKUP_TABLE[92] = 32'h0738A4E1;
      EXP_LOOKUP_TABLE[93] = 32'h06FFC46B;
      EXP_LOOKUP_TABLE[94] = 32'h06C8A3EF;
      EXP_LOOKUP_TABLE[95] = 32'h069335A6;
      EXP_LOOKUP_TABLE[96] = 32'h065F6C33;
      EXP_LOOKUP_TABLE[97] = 32'h062D3AA3;
      EXP_LOOKUP_TABLE[98] = 32'h05FC946A;
      EXP_LOOKUP_TABLE[99] = 32'h05CD6D5F;
      EXP_LOOKUP_TABLE[100] = 32'h059FB9B6;
      EXP_LOOKUP_TABLE[101] = 32'h05736E03;
      EXP_LOOKUP_TABLE[102] = 32'h05487F33;
      EXP_LOOKUP_TABLE[103] = 32'h051EE28A;
      EXP_LOOKUP_TABLE[104] = 32'h04F68DA1;
      EXP_LOOKUP_TABLE[105] = 32'h04CF7661;
      EXP_LOOKUP_TABLE[106] = 32'h04A99306;
      EXP_LOOKUP_TABLE[107] = 32'h0484DA15;
      EXP_LOOKUP_TABLE[108] = 32'h04614261;
      EXP_LOOKUP_TABLE[109] = 32'h043EC303;
      EXP_LOOKUP_TABLE[110] = 32'h041D535C;
      EXP_LOOKUP_TABLE[111] = 32'h03FCEB0F;
      EXP_LOOKUP_TABLE[112] = 32'h03DD8203;
      EXP_LOOKUP_TABLE[113] = 32'h03BF105B;
      EXP_LOOKUP_TABLE[114] = 32'h03A18E7D;
      EXP_LOOKUP_TABLE[115] = 32'h0384F508;
      EXP_LOOKUP_TABLE[116] = 32'h03693CD4;
      EXP_LOOKUP_TABLE[117] = 32'h034E5EF4;
      EXP_LOOKUP_TABLE[118] = 32'h033454B1;
      EXP_LOOKUP_TABLE[119] = 32'h031B1786;
      EXP_LOOKUP_TABLE[120] = 32'h0302A126;
      EXP_LOOKUP_TABLE[121] = 32'h02EAEB72;
      EXP_LOOKUP_TABLE[122] = 32'h02D3F07D;
      EXP_LOOKUP_TABLE[123] = 32'h02BDAA88;
      EXP_LOOKUP_TABLE[124] = 32'h02A81401;
      EXP_LOOKUP_TABLE[125] = 32'h02932782;
      EXP_LOOKUP_TABLE[126] = 32'h027EDFD1;
      EXP_LOOKUP_TABLE[127] = 32'h026B37DB;
      EXP_LOOKUP_TABLE[128] = 32'h02582AB7;
      EXP_LOOKUP_TABLE[129] = 32'h0245B3A0;
      EXP_LOOKUP_TABLE[130] = 32'h0233CDF9;
      EXP_LOOKUP_TABLE[131] = 32'h02227548;
      EXP_LOOKUP_TABLE[132] = 32'h0211A538;
      EXP_LOOKUP_TABLE[133] = 32'h02015994;
      EXP_LOOKUP_TABLE[134] = 32'h01F18E48;
      EXP_LOOKUP_TABLE[135] = 32'h01E23F63;
      EXP_LOOKUP_TABLE[136] = 32'h01D36911;
      EXP_LOOKUP_TABLE[137] = 32'h01C5079B;
      EXP_LOOKUP_TABLE[138] = 32'h01B71769;
      EXP_LOOKUP_TABLE[139] = 32'h01A994FF;
      EXP_LOOKUP_TABLE[140] = 32'h019C7CFD;
      EXP_LOOKUP_TABLE[141] = 32'h018FCC1C;
      EXP_LOOKUP_TABLE[142] = 32'h01837F31;
      EXP_LOOKUP_TABLE[143] = 32'h01779327;
      EXP_LOOKUP_TABLE[144] = 32'h016C0504;
      EXP_LOOKUP_TABLE[145] = 32'h0160D1E4;
      EXP_LOOKUP_TABLE[146] = 32'h0155F6FA;
      EXP_LOOKUP_TABLE[147] = 32'h014B7190;
      EXP_LOOKUP_TABLE[148] = 32'h01413F04;
      EXP_LOOKUP_TABLE[149] = 32'h01375CCA;
      EXP_LOOKUP_TABLE[150] = 32'h012DC868;
      EXP_LOOKUP_TABLE[151] = 32'h01247F7A;
      EXP_LOOKUP_TABLE[152] = 32'h011B7FAD;
      EXP_LOOKUP_TABLE[153] = 32'h0112C6C2;
      EXP_LOOKUP_TABLE[154] = 32'h010A528A;
      EXP_LOOKUP_TABLE[155] = 32'h010220E8;
      EXP_LOOKUP_TABLE[156] = 32'h00FA2FCF;
      EXP_LOOKUP_TABLE[157] = 32'h00F27D44;
      EXP_LOOKUP_TABLE[158] = 32'h00EB075A;
      EXP_LOOKUP_TABLE[159] = 32'h00E3CC32;
      EXP_LOOKUP_TABLE[160] = 32'h00DCC9FF;
      EXP_LOOKUP_TABLE[161] = 32'h00D5FEFF;
      EXP_LOOKUP_TABLE[162] = 32'h00CF6980;
      EXP_LOOKUP_TABLE[163] = 32'h00C907DC;
      EXP_LOOKUP_TABLE[164] = 32'h00C2D87C;
      EXP_LOOKUP_TABLE[165] = 32'h00BCD9D3;
      EXP_LOOKUP_TABLE[166] = 32'h00B70A61;
      EXP_LOOKUP_TABLE[167] = 32'h00B168B3;
      EXP_LOOKUP_TABLE[168] = 32'h00ABF35F;
      EXP_LOOKUP_TABLE[169] = 32'h00A6A90A;
      EXP_LOOKUP_TABLE[170] = 32'h00A18860;
      EXP_LOOKUP_TABLE[171] = 32'h009C9018;
      EXP_LOOKUP_TABLE[172] = 32'h0097BEF6;
      EXP_LOOKUP_TABLE[173] = 32'h009313C4;
      EXP_LOOKUP_TABLE[174] = 32'h008E8D57;
      EXP_LOOKUP_TABLE[175] = 32'h008A2A8F;
      EXP_LOOKUP_TABLE[176] = 32'h0085EA52;
      EXP_LOOKUP_TABLE[177] = 32'h0081CB91;
      EXP_LOOKUP_TABLE[178] = 32'h007DCD43;
      EXP_LOOKUP_TABLE[179] = 32'h0079EE69;
      EXP_LOOKUP_TABLE[180] = 32'h00762E0B;
      EXP_LOOKUP_TABLE[181] = 32'h00728B39;
      EXP_LOOKUP_TABLE[182] = 32'h006F050B;
      EXP_LOOKUP_TABLE[183] = 32'h006B9A9E;
      EXP_LOOKUP_TABLE[184] = 32'h00684B19;
      EXP_LOOKUP_TABLE[185] = 32'h006515A7;
      EXP_LOOKUP_TABLE[186] = 32'h0061F97B;
      EXP_LOOKUP_TABLE[187] = 32'h005EF5CE;
      EXP_LOOKUP_TABLE[188] = 32'h005C09DF;
      EXP_LOOKUP_TABLE[189] = 32'h005934F3;
      EXP_LOOKUP_TABLE[190] = 32'h00567654;
      EXP_LOOKUP_TABLE[191] = 32'h0053CD54;
      EXP_LOOKUP_TABLE[192] = 32'h00513947;
      EXP_LOOKUP_TABLE[193] = 32'h004EB989;
      EXP_LOOKUP_TABLE[194] = 32'h004C4D7A;
      EXP_LOOKUP_TABLE[195] = 32'h0049F47F;
      EXP_LOOKUP_TABLE[196] = 32'h0047AE01;
      EXP_LOOKUP_TABLE[197] = 32'h0045796F;
      EXP_LOOKUP_TABLE[198] = 32'h0043563C;
      EXP_LOOKUP_TABLE[199] = 32'h004143DE;
      EXP_LOOKUP_TABLE[200] = 32'h003F41D2;
      EXP_LOOKUP_TABLE[201] = 32'h003D4F97;
      EXP_LOOKUP_TABLE[202] = 32'h003B6CB0;
      EXP_LOOKUP_TABLE[203] = 32'h003998A4;
      EXP_LOOKUP_TABLE[204] = 32'h0037D2FF;
      EXP_LOOKUP_TABLE[205] = 32'h00361B4F;
      EXP_LOOKUP_TABLE[206] = 32'h00347126;
      EXP_LOOKUP_TABLE[207] = 32'h0032D41A;
      EXP_LOOKUP_TABLE[208] = 32'h003143C3;
      EXP_LOOKUP_TABLE[209] = 32'h002FBFBD;
      EXP_LOOKUP_TABLE[210] = 32'h002E47A7;
      EXP_LOOKUP_TABLE[211] = 32'h002CDB23;
      EXP_LOOKUP_TABLE[212] = 32'h002B79D7;
      EXP_LOOKUP_TABLE[213] = 32'h002A2369;
      EXP_LOOKUP_TABLE[214] = 32'h0028D784;
      EXP_LOOKUP_TABLE[215] = 32'h002795D5;
      EXP_LOOKUP_TABLE[216] = 32'h00265E0C;
      EXP_LOOKUP_TABLE[217] = 32'h00252FDB;
      EXP_LOOKUP_TABLE[218] = 32'h00240AF6;
      EXP_LOOKUP_TABLE[219] = 32'h0022EF14;
      EXP_LOOKUP_TABLE[220] = 32'h0021DBED;
      EXP_LOOKUP_TABLE[221] = 32'h0020D13E;
      EXP_LOOKUP_TABLE[222] = 32'h001FCEC3;
      EXP_LOOKUP_TABLE[223] = 32'h001ED43D;
      EXP_LOOKUP_TABLE[224] = 32'h001DE16B;
      EXP_LOOKUP_TABLE[225] = 32'h001CF612;
      EXP_LOOKUP_TABLE[226] = 32'h001C11F7;
      EXP_LOOKUP_TABLE[227] = 32'h001B34E0;
      EXP_LOOKUP_TABLE[228] = 32'h001A5E96;
      EXP_LOOKUP_TABLE[229] = 32'h00198EE5;
      EXP_LOOKUP_TABLE[230] = 32'h0018C597;
      EXP_LOOKUP_TABLE[231] = 32'h0018027B;
      EXP_LOOKUP_TABLE[232] = 32'h0017455F;
      EXP_LOOKUP_TABLE[233] = 32'h00168E15;
      EXP_LOOKUP_TABLE[234] = 32'h0015DC6F;
      EXP_LOOKUP_TABLE[235] = 32'h00153040;
      EXP_LOOKUP_TABLE[236] = 32'h0014895D;
      EXP_LOOKUP_TABLE[237] = 32'h0013E79C;
      EXP_LOOKUP_TABLE[238] = 32'h00134AD6;
      EXP_LOOKUP_TABLE[239] = 32'h0012B2E2;
      EXP_LOOKUP_TABLE[240] = 32'h00121F9B;
      EXP_LOOKUP_TABLE[241] = 32'h001190DC;
      EXP_LOOKUP_TABLE[242] = 32'h00110682;
      EXP_LOOKUP_TABLE[243] = 32'h00108069;
      EXP_LOOKUP_TABLE[244] = 32'h000FFE70;
      EXP_LOOKUP_TABLE[245] = 32'h000F8077;
      EXP_LOOKUP_TABLE[246] = 32'h000F065E;
      EXP_LOOKUP_TABLE[247] = 32'h000E9007;
      EXP_LOOKUP_TABLE[248] = 32'h000E1D54;
      EXP_LOOKUP_TABLE[249] = 32'h000DAE28;
      EXP_LOOKUP_TABLE[250] = 32'h000D4268;
      EXP_LOOKUP_TABLE[251] = 32'h000CD9F9;
      EXP_LOOKUP_TABLE[252] = 32'h000C74C0;
      EXP_LOOKUP_TABLE[253] = 32'h000C12A5;
      EXP_LOOKUP_TABLE[254] = 32'h000BB38E;
      EXP_LOOKUP_TABLE[255] = 32'h000B5764;
      EXP_LOOKUP_TABLE[256] = 32'h000AFE10;
      EXP_LOOKUP_TABLE[257] = 32'h000AA77C;
      EXP_LOOKUP_TABLE[258] = 32'h000A5391;
      EXP_LOOKUP_TABLE[259] = 32'h000A023C;
      EXP_LOOKUP_TABLE[260] = 32'h0009B367;
      EXP_LOOKUP_TABLE[261] = 32'h000966FF;
      EXP_LOOKUP_TABLE[262] = 32'h00091CF0;
      EXP_LOOKUP_TABLE[263] = 32'h0008D52A;
      EXP_LOOKUP_TABLE[264] = 32'h00088F98;
      EXP_LOOKUP_TABLE[265] = 32'h00084C2A;
      EXP_LOOKUP_TABLE[266] = 32'h00080AD0;
      EXP_LOOKUP_TABLE[267] = 32'h0007CB78;
      EXP_LOOKUP_TABLE[268] = 32'h00078E13;
      EXP_LOOKUP_TABLE[269] = 32'h00075292;
      EXP_LOOKUP_TABLE[270] = 32'h000718E5;
      EXP_LOOKUP_TABLE[271] = 32'h0006E0FF;
      EXP_LOOKUP_TABLE[272] = 32'h0006AAD0;
      EXP_LOOKUP_TABLE[273] = 32'h0006764D;
      EXP_LOOKUP_TABLE[274] = 32'h00064367;
      EXP_LOOKUP_TABLE[275] = 32'h00061212;
      EXP_LOOKUP_TABLE[276] = 32'h0005E242;
      EXP_LOOKUP_TABLE[277] = 32'h0005B3EA;
      EXP_LOOKUP_TABLE[278] = 32'h00058700;
      EXP_LOOKUP_TABLE[279] = 32'h00055B77;
      EXP_LOOKUP_TABLE[280] = 32'h00053145;
      EXP_LOOKUP_TABLE[281] = 32'h0005085F;
      EXP_LOOKUP_TABLE[282] = 32'h0004E0BB;
      EXP_LOOKUP_TABLE[283] = 32'h0004BA50;
      EXP_LOOKUP_TABLE[284] = 32'h00049513;
      EXP_LOOKUP_TABLE[285] = 32'h000470FC;
      EXP_LOOKUP_TABLE[286] = 32'h00044E00;
      EXP_LOOKUP_TABLE[287] = 32'h00042C19;
      EXP_LOOKUP_TABLE[288] = 32'h00040B3C;
      EXP_LOOKUP_TABLE[289] = 32'h0003EB62;
      EXP_LOOKUP_TABLE[290] = 32'h0003CC83;
      EXP_LOOKUP_TABLE[291] = 32'h0003AE97;
      EXP_LOOKUP_TABLE[292] = 32'h00039197;
      EXP_LOOKUP_TABLE[293] = 32'h0003757C;
      EXP_LOOKUP_TABLE[294] = 32'h00035A3D;
      EXP_LOOKUP_TABLE[295] = 32'h00033FD5;
      EXP_LOOKUP_TABLE[296] = 32'h0003263E;
      EXP_LOOKUP_TABLE[297] = 32'h00030D6F;
      EXP_LOOKUP_TABLE[298] = 32'h0002F565;
      EXP_LOOKUP_TABLE[299] = 32'h0002DE17;
      EXP_LOOKUP_TABLE[300] = 32'h0002C781;
      EXP_LOOKUP_TABLE[301] = 32'h0002B19D;
      EXP_LOOKUP_TABLE[302] = 32'h00029C66;
      EXP_LOOKUP_TABLE[303] = 32'h000287D5;
      EXP_LOOKUP_TABLE[304] = 32'h000273E7;
      EXP_LOOKUP_TABLE[305] = 32'h00026095;
      EXP_LOOKUP_TABLE[306] = 32'h00024DDC;
      EXP_LOOKUP_TABLE[307] = 32'h00023BB6;
      EXP_LOOKUP_TABLE[308] = 32'h00022A1F;
      EXP_LOOKUP_TABLE[309] = 32'h00021912;
      EXP_LOOKUP_TABLE[310] = 32'h0002088C;
      EXP_LOOKUP_TABLE[311] = 32'h0001F888;
      EXP_LOOKUP_TABLE[312] = 32'h0001E902;
      EXP_LOOKUP_TABLE[313] = 32'h0001D9F7;
      EXP_LOOKUP_TABLE[314] = 32'h0001CB62;
      EXP_LOOKUP_TABLE[315] = 32'h0001BD3F;
      EXP_LOOKUP_TABLE[316] = 32'h0001AF8C;
      EXP_LOOKUP_TABLE[317] = 32'h0001A245;
      EXP_LOOKUP_TABLE[318] = 32'h00019567;
      EXP_LOOKUP_TABLE[319] = 32'h000188EE;
      EXP_LOOKUP_TABLE[320] = 32'h00017CD7;
      EXP_LOOKUP_TABLE[321] = 32'h0001711F;
      EXP_LOOKUP_TABLE[322] = 32'h000165C4;
      EXP_LOOKUP_TABLE[323] = 32'h00015AC2;
      EXP_LOOKUP_TABLE[324] = 32'h00015017;
      EXP_LOOKUP_TABLE[325] = 32'h000145C0;
      EXP_LOOKUP_TABLE[326] = 32'h00013BBA;
      EXP_LOOKUP_TABLE[327] = 32'h00013203;
      EXP_LOOKUP_TABLE[328] = 32'h00012899;
      EXP_LOOKUP_TABLE[329] = 32'h00011F79;
      EXP_LOOKUP_TABLE[330] = 32'h000116A1;
      EXP_LOOKUP_TABLE[331] = 32'h00010E0E;
      EXP_LOOKUP_TABLE[332] = 32'h000105BF;
      EXP_LOOKUP_TABLE[333] = 32'h0000FDB2;
      EXP_LOOKUP_TABLE[334] = 32'h0000F5E3;
      EXP_LOOKUP_TABLE[335] = 32'h0000EE53;
      EXP_LOOKUP_TABLE[336] = 32'h0000E6FE;
      EXP_LOOKUP_TABLE[337] = 32'h0000DFE2;
      EXP_LOOKUP_TABLE[338] = 32'h0000D8FF;
      EXP_LOOKUP_TABLE[339] = 32'h0000D252;
      EXP_LOOKUP_TABLE[340] = 32'h0000CBD9;
      EXP_LOOKUP_TABLE[341] = 32'h0000C594;
      EXP_LOOKUP_TABLE[342] = 32'h0000BF7F;
      EXP_LOOKUP_TABLE[343] = 32'h0000B99B;
      EXP_LOOKUP_TABLE[344] = 32'h0000B3E5;
      EXP_LOOKUP_TABLE[345] = 32'h0000AE5C;
      EXP_LOOKUP_TABLE[346] = 32'h0000A8FF;
      EXP_LOOKUP_TABLE[347] = 32'h0000A3CC;
      EXP_LOOKUP_TABLE[348] = 32'h00009EC2;
      EXP_LOOKUP_TABLE[349] = 32'h000099DF;
      EXP_LOOKUP_TABLE[350] = 32'h00009523;
      EXP_LOOKUP_TABLE[351] = 32'h0000908D;
      EXP_LOOKUP_TABLE[352] = 32'h00008C1A;
      EXP_LOOKUP_TABLE[353] = 32'h000087CB;
      EXP_LOOKUP_TABLE[354] = 32'h0000839D;
      EXP_LOOKUP_TABLE[355] = 32'h00007F90;
      EXP_LOOKUP_TABLE[356] = 32'h00007BA4;
      EXP_LOOKUP_TABLE[357] = 32'h000077D6;
      EXP_LOOKUP_TABLE[358] = 32'h00007426;
      EXP_LOOKUP_TABLE[359] = 32'h00007093;
      EXP_LOOKUP_TABLE[360] = 32'h00006D1C;
      EXP_LOOKUP_TABLE[361] = 32'h000069C1;
      EXP_LOOKUP_TABLE[362] = 32'h00006680;
      EXP_LOOKUP_TABLE[363] = 32'h00006359;
      EXP_LOOKUP_TABLE[364] = 32'h0000604A;
      EXP_LOOKUP_TABLE[365] = 32'h00005D54;
      EXP_LOOKUP_TABLE[366] = 32'h00005A75;
      EXP_LOOKUP_TABLE[367] = 32'h000057AC;
      EXP_LOOKUP_TABLE[368] = 32'h000054FA;
      EXP_LOOKUP_TABLE[369] = 32'h0000525C;
      EXP_LOOKUP_TABLE[370] = 32'h00004FD4;
      EXP_LOOKUP_TABLE[371] = 32'h00004D5F;
      EXP_LOOKUP_TABLE[372] = 32'h00004AFE;
      EXP_LOOKUP_TABLE[373] = 32'h000048AF;
      EXP_LOOKUP_TABLE[374] = 32'h00004672;
      EXP_LOOKUP_TABLE[375] = 32'h00004447;
      EXP_LOOKUP_TABLE[376] = 32'h0000422E;
      EXP_LOOKUP_TABLE[377] = 32'h00004024;
      EXP_LOOKUP_TABLE[378] = 32'h00003E2B;
      EXP_LOOKUP_TABLE[379] = 32'h00003C42;
      EXP_LOOKUP_TABLE[380] = 32'h00003A67;
      EXP_LOOKUP_TABLE[381] = 32'h0000389B;
      EXP_LOOKUP_TABLE[382] = 32'h000036DD;
      EXP_LOOKUP_TABLE[383] = 32'h0000352D;
      EXP_LOOKUP_TABLE[384] = 32'h0000338A;
      EXP_LOOKUP_TABLE[385] = 32'h000031F4;
      EXP_LOOKUP_TABLE[386] = 32'h0000306B;
      EXP_LOOKUP_TABLE[387] = 32'h00002EED;
      EXP_LOOKUP_TABLE[388] = 32'h00002D7C;
      EXP_LOOKUP_TABLE[389] = 32'h00002C15;
      EXP_LOOKUP_TABLE[390] = 32'h00002ABA;
      EXP_LOOKUP_TABLE[391] = 32'h0000296A;
      EXP_LOOKUP_TABLE[392] = 32'h00002823;
      EXP_LOOKUP_TABLE[393] = 32'h000026E7;
      EXP_LOOKUP_TABLE[394] = 32'h000025B5;
      EXP_LOOKUP_TABLE[395] = 32'h0000248C;
      EXP_LOOKUP_TABLE[396] = 32'h0000236C;
      EXP_LOOKUP_TABLE[397] = 32'h00002255;
      EXP_LOOKUP_TABLE[398] = 32'h00002147;
      EXP_LOOKUP_TABLE[399] = 32'h00002040;
      EXP_LOOKUP_TABLE[400] = 32'h00001F42;
      EXP_LOOKUP_TABLE[401] = 32'h00001E4C;
      EXP_LOOKUP_TABLE[402] = 32'h00001D5E;
      EXP_LOOKUP_TABLE[403] = 32'h00001C76;
      EXP_LOOKUP_TABLE[404] = 32'h00001B96;
      EXP_LOOKUP_TABLE[405] = 32'h00001ABD;
      EXP_LOOKUP_TABLE[406] = 32'h000019EA;
      EXP_LOOKUP_TABLE[407] = 32'h0000191E;
      EXP_LOOKUP_TABLE[408] = 32'h00001858;
      EXP_LOOKUP_TABLE[409] = 32'h00001798;
      EXP_LOOKUP_TABLE[410] = 32'h000016DF;
      EXP_LOOKUP_TABLE[411] = 32'h0000162A;
      EXP_LOOKUP_TABLE[412] = 32'h0000157C;
      EXP_LOOKUP_TABLE[413] = 32'h000014D3;
      EXP_LOOKUP_TABLE[414] = 32'h0000142F;
      EXP_LOOKUP_TABLE[415] = 32'h00001390;
      EXP_LOOKUP_TABLE[416] = 32'h000012F6;
      EXP_LOOKUP_TABLE[417] = 32'h00001260;
      EXP_LOOKUP_TABLE[418] = 32'h000011CF;
      EXP_LOOKUP_TABLE[419] = 32'h00001143;
      EXP_LOOKUP_TABLE[420] = 32'h000010BB;
      EXP_LOOKUP_TABLE[421] = 32'h00001037;
      EXP_LOOKUP_TABLE[422] = 32'h00000FB8;
      EXP_LOOKUP_TABLE[423] = 32'h00000F3C;
      EXP_LOOKUP_TABLE[424] = 32'h00000EC4;
      EXP_LOOKUP_TABLE[425] = 32'h00000E50;
      EXP_LOOKUP_TABLE[426] = 32'h00000DDF;
      EXP_LOOKUP_TABLE[427] = 32'h00000D72;
      EXP_LOOKUP_TABLE[428] = 32'h00000D08;
      EXP_LOOKUP_TABLE[429] = 32'h00000CA1;
      EXP_LOOKUP_TABLE[430] = 32'h00000C3D;
      EXP_LOOKUP_TABLE[431] = 32'h00000BDD;
      EXP_LOOKUP_TABLE[432] = 32'h00000B80;
      EXP_LOOKUP_TABLE[433] = 32'h00000B25;
      EXP_LOOKUP_TABLE[434] = 32'h00000ACD;
      EXP_LOOKUP_TABLE[435] = 32'h00000A78;
      EXP_LOOKUP_TABLE[436] = 32'h00000A26;
      EXP_LOOKUP_TABLE[437] = 32'h000009D6;
      EXP_LOOKUP_TABLE[438] = 32'h00000988;
      EXP_LOOKUP_TABLE[439] = 32'h0000093D;
      EXP_LOOKUP_TABLE[440] = 32'h000008F4;
      EXP_LOOKUP_TABLE[441] = 32'h000008AE;
      EXP_LOOKUP_TABLE[442] = 32'h00000869;
      EXP_LOOKUP_TABLE[443] = 32'h00000827;
      EXP_LOOKUP_TABLE[444] = 32'h000007E7;
      EXP_LOOKUP_TABLE[445] = 32'h000007A9;
      EXP_LOOKUP_TABLE[446] = 32'h0000076C;
      EXP_LOOKUP_TABLE[447] = 32'h00000732;
      EXP_LOOKUP_TABLE[448] = 32'h000006F9;
      EXP_LOOKUP_TABLE[449] = 32'h000006C2;
      EXP_LOOKUP_TABLE[450] = 32'h0000068D;
      EXP_LOOKUP_TABLE[451] = 32'h00000659;
      EXP_LOOKUP_TABLE[452] = 32'h00000627;
      EXP_LOOKUP_TABLE[453] = 32'h000005F7;
      EXP_LOOKUP_TABLE[454] = 32'h000005C8;
      EXP_LOOKUP_TABLE[455] = 32'h0000059A;
      EXP_LOOKUP_TABLE[456] = 32'h0000056E;
      EXP_LOOKUP_TABLE[457] = 32'h00000543;
      EXP_LOOKUP_TABLE[458] = 32'h0000051A;
      EXP_LOOKUP_TABLE[459] = 32'h000004F2;
      EXP_LOOKUP_TABLE[460] = 32'h000004CB;
      EXP_LOOKUP_TABLE[461] = 32'h000004A5;
      EXP_LOOKUP_TABLE[462] = 32'h00000480;
      EXP_LOOKUP_TABLE[463] = 32'h0000045D;
      EXP_LOOKUP_TABLE[464] = 32'h0000043B;
      EXP_LOOKUP_TABLE[465] = 32'h00000419;
      EXP_LOOKUP_TABLE[466] = 32'h000003F9;
      EXP_LOOKUP_TABLE[467] = 32'h000003DA;
      EXP_LOOKUP_TABLE[468] = 32'h000003BB;
      EXP_LOOKUP_TABLE[469] = 32'h0000039E;
      EXP_LOOKUP_TABLE[470] = 32'h00000381;
      EXP_LOOKUP_TABLE[471] = 32'h00000366;
      EXP_LOOKUP_TABLE[472] = 32'h0000034B;
      EXP_LOOKUP_TABLE[473] = 32'h00000331;
      EXP_LOOKUP_TABLE[474] = 32'h00000318;
      EXP_LOOKUP_TABLE[475] = 32'h00000300;
      EXP_LOOKUP_TABLE[476] = 32'h000002E8;
      EXP_LOOKUP_TABLE[477] = 32'h000002D1;
      EXP_LOOKUP_TABLE[478] = 32'h000002BB;
      EXP_LOOKUP_TABLE[479] = 32'h000002A5;
      EXP_LOOKUP_TABLE[480] = 32'h00000290;
      EXP_LOOKUP_TABLE[481] = 32'h0000027C;
      EXP_LOOKUP_TABLE[482] = 32'h00000269;
      EXP_LOOKUP_TABLE[483] = 32'h00000256;
      EXP_LOOKUP_TABLE[484] = 32'h00000243;
      EXP_LOOKUP_TABLE[485] = 32'h00000231;
      EXP_LOOKUP_TABLE[486] = 32'h00000220;
      EXP_LOOKUP_TABLE[487] = 32'h0000020F;
      EXP_LOOKUP_TABLE[488] = 32'h000001FF;
      EXP_LOOKUP_TABLE[489] = 32'h000001EF;
      EXP_LOOKUP_TABLE[490] = 32'h000001E0;
      EXP_LOOKUP_TABLE[491] = 32'h000001D1;
      EXP_LOOKUP_TABLE[492] = 32'h000001C3;
      EXP_LOOKUP_TABLE[493] = 32'h000001B5;
      EXP_LOOKUP_TABLE[494] = 32'h000001A8;
      EXP_LOOKUP_TABLE[495] = 32'h0000019B;
      EXP_LOOKUP_TABLE[496] = 32'h0000018E;
      EXP_LOOKUP_TABLE[497] = 32'h00000182;
      EXP_LOOKUP_TABLE[498] = 32'h00000176;
      EXP_LOOKUP_TABLE[499] = 32'h0000016A;
      EXP_LOOKUP_TABLE[500] = 32'h0000015F;
      EXP_LOOKUP_TABLE[501] = 32'h00000154;
      EXP_LOOKUP_TABLE[502] = 32'h0000014A;
      EXP_LOOKUP_TABLE[503] = 32'h00000140;
      EXP_LOOKUP_TABLE[504] = 32'h00000136;
      EXP_LOOKUP_TABLE[505] = 32'h0000012C;
      EXP_LOOKUP_TABLE[506] = 32'h00000123;
      EXP_LOOKUP_TABLE[507] = 32'h0000011A;
      EXP_LOOKUP_TABLE[508] = 32'h00000111;
      EXP_LOOKUP_TABLE[509] = 32'h00000109;
      EXP_LOOKUP_TABLE[510] = 32'h00000101;
      EXP_LOOKUP_TABLE[511] = 32'h000000F9;
      EXP_LOOKUP_TABLE[512] = 32'h000000F1;
  end

  wire [31:0] frac_bits = cmd_payload_inputs_0;
  wire [31:0] raw_input = cmd_payload_inputs_1;

  parameter [1:0] EXP_in = 2'b00;

  wire [31:0] exp_index;
  parameter [12:0] exp_table_size = 512;  // 2^9
  parameter [4:0] exp_table_offset_bit = 5;  // 因為輸入絕對值範圍為 0~16，所以offset bit設為 9 - 4 = 5

  assign exp_index = (~raw_input + 1) >> (frac_bits - exp_table_offset_bit);
  
   // Only not ready for a command when we have a response.
  assign cmd_ready = ~rsp_valid;

  always @(posedge clk) begin
    if (reset) begin
      rsp_payload_outputs_0 <= 0;
      rsp_valid <= 0;
    end else if (rsp_valid) begin
      rsp_valid <= ~rsp_ready;
    end else if (cmd_valid) begin
      rsp_valid <= 1;
      case (cmd_payload_function_id[9:3])
        EXP_in: begin
          rsp_payload_outputs_0 <= EXP_LOOKUP_TABLE[(exp_index < exp_table_size) ? exp_index : exp_table_size - 1];
        end
        default: begin
        end
      endcase
    end
  end

endmodule
